// `defines are written for the asynchronous fifo

`define DATA_WIDTH 8